module T_flipflop (
 input clk, rst_n,
 input t,
 output reg q,
 output q_bar
 );
 
 // always@(posedge clk or negedge rst_n) // for asynchronous reset
 always@(posedge clk) begin // for synchronous reset
 if(!rst_n) q <= 0;
 else begin
 q <= (t?~q:q);
 end
 end
 assign q_bar = ~q;
endmodule
